Name,SN,Age,Address
Chor,1,23,Kathmandu
Shyam,2,45,Bara
Nabin,3,54,Pokhara
Santosh,4,45,Slolu
